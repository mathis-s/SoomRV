module ReservationStation
#(
    parameter QUEUE_SIZE = 1;
)
(
    input wire clk,
    input wire rst,

    input UOp uop,
    
);