`include "src/Include.sv"

module Rename
(
    
);



endmodule