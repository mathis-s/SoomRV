module IssueQueue
#(
    parameter SIZE = 8,
    parameter NUM_OPERANDS = 2,
    parameter NUM_UOPS = 4,
    parameter RESULT_BUS_COUNT = 4,
    parameter IMM_BITS=32,
    parameter FU0 = FU_ST,
    parameter FU1 = FU_ST,
    parameter FU2 = FU_ST,
    parameter FU3 = FU_ST,
    parameter FU0_SPLIT=0,
    parameter FU0_ORDER=0,
    parameter FU1_DLY=0
    
)
(
    input wire clk,
    input wire rst,
    input wire frontEn,
    
    input wire IN_stall,
    input wire IN_doNotIssueFU1,
    input wire IN_doNotIssueFU2,
    
    input wire IN_uopValid[NUM_UOPS-1:0],
    input R_UOp IN_uop[NUM_UOPS-1:0],
    input wire IN_uopOrdering[NUM_UOPS-1:0],
    
    input wire IN_resultValid[RESULT_BUS_COUNT-1:0],
    input RES_UOp IN_resultUOp[RESULT_BUS_COUNT-1:0],
    
    input wire IN_loadForwardValid,
    input Tag IN_loadForwardTag,
    
    input BranchProv IN_branch,
    
    // All ops that are being issued (including OUT_uop)
    // For operand forwarding
    input wire IN_issueValid[NUM_UOPS-1:0],
    input R_UOp IN_issueUOps[NUM_UOPS-1:0],
    
    input SqN IN_maxStoreSqN,
    input SqN IN_maxLoadSqN,
    
    output reg OUT_valid,
    output R_UOp OUT_uop,
    
    output reg OUT_full
);

localparam ID_LEN = $clog2(SIZE);

integer i;
integer j;
integer k;

typedef struct packed
{
    logic[IMM_BITS-1:0] imm;
    
    logic[NUM_OPERANDS-1:0] avail;
    Tag[NUM_OPERANDS-1:0] tags;
    
    logic immB;
    SqN sqN;
    Tag tagDst;
    RegNm nmDst;
    logic[5:0] opcode;
    FetchID_t fetchID;
    FetchOff_t fetchOffs;
    SqN storeSqN;
    SqN loadSqN;
    FuncUnit fu;
    logic compressed;
} R_ST_UOp;

R_ST_UOp queue[SIZE-1:0];
reg valid[SIZE-1:0];

reg[$clog2(SIZE):0] insertIndex;
reg[32:0] reservedWBs;

//assign OUT_full = insertIndex > (SIZE-NUM_UOPS);

reg[NUM_OPERANDS-1:0] newAvail[SIZE-1:0];
reg[NUM_OPERANDS-1:0] newAvail_dl[SIZE-1:0];


always_comb begin
    for (i = 0; i < SIZE; i=i+1) begin
        
        for (k = 0; k < NUM_OPERANDS; k=k+1) begin
            newAvail[i][k] = 0;
            newAvail_dl[i][k] = 0;
        end
        
        for (j = 0; j < RESULT_BUS_COUNT; j=j+1) begin
            for (k = 0; k < NUM_OPERANDS; k=k+1)
                if (IN_resultValid[j] && queue[i].tags[k] == IN_resultUOp[j].tagDst) newAvail[i][k] = 1;
        end
        
        for (j = 0; j < 2; j=j+1) begin
            if (IN_issueValid[j] && IN_issueUOps[j].nmDst != 0) begin
                if (IN_issueUOps[j].fu == FU_INT) begin
                    for (k = 0; k < NUM_OPERANDS; k=k+1)
                        if (queue[i].tags[k] == IN_issueUOps[j].tagDst) newAvail[i][k] = 1;
                end
                else if (IN_issueUOps[j].fu == FU_FPU || IN_issueUOps[j].fu == FU_FMUL) begin
                    for (k = 0; k < NUM_OPERANDS; k=k+1)
                        if (queue[i].tags[k] == IN_issueUOps[j].tagDst) newAvail_dl[i][k] = 1;
                end
            end
        end
        
        for (k = 0; k < NUM_OPERANDS; k=k+1)
            if (IN_loadForwardValid && queue[i].tags[k] == IN_loadForwardTag) newAvail[i][k] = 1;
    end
end

always_comb begin
    reg[$clog2(SIZE):0] count = 0;
    for (i = 0; i < NUM_UOPS; i=i+1) begin
        if (IN_uopValid[i] && 
            ((IN_uop[i].fu == FU0 && (!FU0_SPLIT || IN_uopOrdering[i] == FU0_ORDER)) || 
                IN_uop[i].fu == FU1 || IN_uop[i].fu == FU2 || IN_uop[i].fu == FU3)) begin
            count = count + 1;
        end
    end
    OUT_full = insertIndex > (SIZE[$clog2(SIZE):0] - count);
end

always_ff@(posedge clk) begin
    
    // Update availability
    for (i = 0; i < SIZE; i=i+1) begin
        queue[i].avail <= queue[i].avail | newAvail[i] | newAvail_dl[i];
    end
    reservedWBs <= {1'b0, reservedWBs[32:1]};
    
    if (rst) begin
        insertIndex = 0;
        reservedWBs <= 0;
        OUT_valid <= 0;
    end
    else if (IN_branch.taken) begin
        
        reg[ID_LEN:0] newInsertIndex = 0;
        // Set insert index to first invalid entry
        for (i = 0; i < SIZE; i=i+1) begin
            if (i < insertIndex && $signed(queue[i].sqN - IN_branch.sqN) <= 0) begin
                newInsertIndex = i[$clog2(SIZE):0] + 1;
            end
        end
        insertIndex = newInsertIndex;
        if (!IN_stall || $signed(OUT_uop.sqN - IN_branch.sqN) > 0)
            OUT_valid <= 0;
    end
    else begin
        reg issued = 0;
        
        // Issue
        if (!IN_stall) begin
            OUT_valid <= 0;
            
            for (i = 0; i < SIZE; i=i+1) begin
                if (i < insertIndex && !issued) begin
                    if (&(queue[i].avail | newAvail[i]) &&
                        (queue[i].fu != FU1 || !IN_doNotIssueFU1) && 
                        (queue[i].fu != FU2 || !IN_doNotIssueFU2) && 
                        !((queue[i].fu == FU_INT || queue[i].fu == FU_FPU || queue[i].fu == FU_FMUL) && reservedWBs[0]) && 
                        
                        // Only issue stores that fit into store queue
                        ((FU0 != FU_ST && FU1 != FU_ST && FU2 != FU_ST && FU3 != FU_ST) || 
                            queue[i].fu != FU_ST || $signed(queue[i].storeSqN - IN_maxStoreSqN) <= 0) &&
                        
                        // Only issue loads that fit into load order buffer
                        ((FU0 != FU_LD && FU1 != FU_LD && FU2 != FU_LD && FU3 != FU_LD) || 
                            queue[i].fu != FU_LD || $signed(queue[i].loadSqN - IN_maxLoadSqN) <= 0)) begin
                        
                        issued = 1;
                        OUT_valid <= 1;
                        //OUT_uop <= queue[i];
                        
                        OUT_uop.imm <= {{(32 - IMM_BITS){1'b0}}, queue[i].imm};
                        
                        OUT_uop.availA <= queue[i].avail[0];
                        OUT_uop.tagA <= queue[i].tags[0];
                        
                        if (NUM_OPERANDS >= 2) begin
                            // verilator lint_off SELRANGE
                            OUT_uop.availB <= queue[i].avail[1];
                            OUT_uop.tagB <= queue[i].tags[1];
                            // verilator lint_on SELRANGE
                        end
                        else begin
                            OUT_uop.availB <= 1;
                            OUT_uop.tagB <= 7'h40;
                        end
                        
                        OUT_uop.immB <= queue[i].immB;
                        OUT_uop.sqN <= queue[i].sqN;
                        OUT_uop.tagDst <= queue[i].tagDst;
                        OUT_uop.nmDst <= queue[i].nmDst;
                        OUT_uop.opcode <= queue[i].opcode;
                        OUT_uop.fetchID <= queue[i].fetchID;
                        OUT_uop.fetchOffs <= queue[i].fetchOffs;
                        OUT_uop.storeSqN <= queue[i].storeSqN;
                        OUT_uop.loadSqN <= queue[i].loadSqN;
                        OUT_uop.fu <= queue[i].fu;
                        OUT_uop.compressed <= queue[i].compressed;
                        
                        // Shift other ops forward
                        for (j = i; j < SIZE-1; j=j+1) begin
                            queue[j] <= queue[j+1];
                            queue[j].avail <= queue[j+1].avail | newAvail[j+1] | newAvail_dl[j+1];
                        end
                        insertIndex = insertIndex - 1;
                        
                        // Reserve WB if this is a slow operation
                        if (queue[i].fu == FU1 && FU1_DLY > 0)
                            reservedWBs <= {1'b0, reservedWBs[32:1]} | (1 << (FU1_DLY - 1));
                    end
                end
            end
        end
        
        // Enqueue
        if (frontEn) begin
            for (i = 0; i < NUM_UOPS; i=i+1) begin
                if (IN_uopValid[i] && 
                    ((IN_uop[i].fu == FU0 && (!FU0_SPLIT || IN_uopOrdering[i] == FU0_ORDER)) || 
                        IN_uop[i].fu == FU1 || IN_uop[i].fu == FU2 || IN_uop[i].fu == FU3)) begin
                    
                    R_ST_UOp temp;// = IN_uop[i];
                    
                    temp.imm = IN_uop[i].imm[IMM_BITS-1:0];
                    
                    temp.avail[0] = IN_uop[i].availA;
                    temp.tags[0] = IN_uop[i].tagA;
                    
                    if (NUM_OPERANDS >= 2) begin
                        // verilator lint_off SELRANGE
                        temp.avail[1] = IN_uop[i].availB;
                        temp.tags[1] = IN_uop[i].tagB;
                        // verilator lint_on SELRANGE
                    end
                    
                    temp.immB = IN_uop[i].immB;
                    temp.sqN = IN_uop[i].sqN;
                    temp.tagDst = IN_uop[i].tagDst;
                    temp.nmDst = IN_uop[i].nmDst;
                    temp.opcode = IN_uop[i].opcode;
                    temp.fetchID = IN_uop[i].fetchID;
                    temp.fetchOffs = IN_uop[i].fetchOffs;
                    temp.storeSqN = IN_uop[i].storeSqN;
                    temp.loadSqN = IN_uop[i].loadSqN;
                    temp.fu = IN_uop[i].fu;
                    temp.compressed = IN_uop[i].compressed;
                    
                    
                    // Check if the result for this op is being broadcasted in the current cycle
                    for (j = 0; j < RESULT_BUS_COUNT; j=j+1) begin
                        if (IN_resultValid[j]) begin
                            for (k = 0; k < NUM_OPERANDS; k=k+1)
                                if (temp.tags[k] == IN_resultUOp[j].tagDst) temp.avail[k] = 1;
                        end
                    end
                    
                    // Special handling for multi-uop instructions
                    if (IN_uop[i].fu == FU_ATOMIC) begin
                    
                        // First uop goes into load FU
                        if (FU0 == FU_LD) begin
                            // Operand is not required
                            // verilator lint_off SELRANGE
                            // temp.tags[1] = 7'h40;
                            // temp.avail[1] = 1;
                            // verilator lint_on SELRANGE
                        end
                        
                        // Second uop goes into first int FU
                        /*else if (FU0 == FU_INT) begin
                            // First operand is loaded value
                            temp.tagA = IN_uop[i].tagDst;
                        end*/
                        
                        // Third uop goes into store FU
                        else if (FU0 == FU_ST) begin
                            // Data operand is result of op
                            //temp.tagB = IN_uop[i].tagDst;
                            //temp.availB = 0;
                            // Result was already written by second uop
                            temp.nmDst = 0;
                        end
                    end
                    
                    queue[insertIndex[ID_LEN-1:0]] <= temp;
                    
                    insertIndex = insertIndex + 1;
                end
            end
        end
    end
end

endmodule
