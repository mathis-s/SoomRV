module RF
(
    
);


endmodule