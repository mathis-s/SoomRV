module Rename
(
    
);



endmodule